LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY mux IS
	PORT(E0, E1, E2, E3, E4, E5, E6, E7, E8 :IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		MC : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END mux;

ARCHITECTURE Behavior OF mux IS

BEGIN
	
		S <= "00000000" WHEN MC = "000000000" ELSE
				E0 WHEN MC = "100000000" ELSE
				E1 WHEN MC = "010000000" ELSE
				E2 WHEN MC = "001000000" ELSE
				E3 WHEN MC = "000100000" ELSE
				E4 WHEN MC = "000010000" ELSE
				E5 WHEN MC = "000001000" ELSE
				E6 WHEN MC = "000000100" ELSE
				E7 WHEN MC = "000000010" ELSE
				E8 WHEN MC = "000000001";
				
END Behavior;