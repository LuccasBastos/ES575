LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY display IS
	PORT(S :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		H: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END display;

ARCHITECTURE Behavior OF display IS

BEGIN
	
	H <= "1000000" WHEN S = "0000" ELSE
				"1111001" WHEN S = "0001" ELSE
				"0100100" WHEN S = "0010" ELSE
				"0110000" WHEN S = "0011" ELSE
				"0011001" WHEN S = "0100" ELSE
				"0010010" WHEN S = "0101" ELSE
				"0000010" WHEN S = "0110" ELSE
				"1111000" WHEN S = "0111" ELSE
				"0000000" WHEN S = "1000" ELSE
				"0010000" WHEN S = "1001" ELSE
				"0001000" WHEN S = "1010" ELSE
				"0000011" WHEN S = "1011" ELSE
				"0100111" WHEN S = "1100" ELSE
				"0100001" WHEN S = "1101" ELSE
				"0000110" WHEN S = "1110" ELSE
				"0001110";
					

END Behavior;